* MAX4040 MACRO MODEL, SINGLE-POLE 
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   vcc
*                   |   |   |	vee
*		    |   |   |   |   output
*		    |   |   |   |   |
.SUBCKT MAX4040	    1   2   0	0   6
* INPUT IMPEDANCE
RIN	1	2	44k
* DC GAIN=20K AND POLE1=4.5Hz
* UNITY GAIN = DCGAIN X POLE1 = 90kHz
EGAIN	3 0	1 2	20k
RP1	3	4	1K
CP1	4	0	35.4uF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER	5 0	4 0	1
ROUT	5	6	100
.ENDS

